// Hello World - Example
module hello_world();

  // Displays the message in the console on a new line with a TAB before
  initial begin
    $display(("\n\t Hello world! \n");
	
  end

endmodule
